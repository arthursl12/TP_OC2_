`ifndef MEM_ONE
`define MEM_ONE

`include "./src/MemoryModule.v"

module Mem_1 (
    input clock,
    input reset,
    input mem_ram_load,

    input m0_m1_oper,
    input m0_m1_readmem,
    input m0_m1_writemem,
    input [31:0] m0_m1_data_addr,
    input [31:0] m0_m1_regb,
    input [4:0] m0_m1_regdest,
    input m0_m1_writereg,

    output reg m1_m2_oper,
    output reg [4:0] m1_m2_regdest,
    output reg m1_m2_writereg,
    output reg [31:0] m1_m2_wbvalue
);

    wire [6:0] data_addr;
    assign data_addr = m0_m1_data_addr[8:2];

    wire data_wre;
    // WRITE flag to memory module
    assign data_wre = !m0_m1_readmem & m0_m1_writemem;

    wire [31:0] data_data_out;

    MemoryModule data_memory (
        .clk(clock),
        .addr(data_addr),
        .data(data_data_out),
        .data_in(m0_m1_regb),
        .write_enable(data_wre)
    );

    // Ram data_ram (
    //     .clock(clock),
    //     .reset(reset),
    //     .addr(data_addr),
    //     .data_in(m0_m1_regb),
    //     .data_out(data_data_out),
    //     .wre(data_wre),
    //     .instr_load(1'b0),
    //     .data_load(mem_ram_load)
    // );

    always @(posedge clock or negedge reset) begin
        if (~reset) begin
            m1_m2_oper <= 1'b0;
            m1_m2_regdest <= 5'b00000;
            m1_m2_writereg <= 1'b0;
            m1_m2_wbvalue <= 32'h0000_0000;
        end else if (~m0_m1_oper) begin
            m1_m2_oper <= 1'b0;
            m1_m2_regdest <= 5'b00000;
            m1_m2_writereg <= 1'b0;
            m1_m2_wbvalue <= 32'h0000_0000;
        end else begin
            m1_m2_oper <= 1'b1;
            m1_m2_regdest <= m0_m1_regdest;
            m1_m2_writereg <= m0_m1_writereg;
            m1_m2_wbvalue <= data_data_out;
        end
    end
   
endmodule

`endif
